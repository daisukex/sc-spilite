class ahbm_agent extends uvm_agent;
  `uvm_component_utils(ahbm_agent)

  function new (string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
  endfunction

endclass
