`include "ahbm_agent.sv"
